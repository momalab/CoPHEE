/**********************************************************************************
    This module is part of the project CoPHEE.
    CoPHEE: A co-processor for partially homomorphic encrypted encryption
    Copyright (C) 2019  Michail Maniatakos
    New York University Abu Dhabi, wp.nyu.edu/momalab/

    If find any of our work useful, please cite our publication:
      M. Nabeel, M. Ashraf, E. Chielle, N.G. Tsoutsos, and M. Maniatakos.
      "CoPHEE: Co-processor for Partially Homomorphic Encrypted Execution". 
      In: IEEE Hardware-Oriented Security and Trust (HOST). 

    This program is free software: you can redistribute it and/or modify
    it under the terms of the GNU General Public License as published by
    the Free Software Foundation, either version 3 of the License, or
    (at your option) any later version.

    This program is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public License for more details.

    You should have received a copy of the GNU General Public License
    along with this program.  If not, see <http://www.gnu.org/licenses/>.
**********************************************************************************/


parameter GPCFG0_ADDR   = 16'h0000;  //PAD03_CTL  UARTM_TX  0_0001_0000
  parameter GPCFG1_ADDR   = 16'h0004;  //PAD04_CTL  UARTM_RX  0_0000_0111
  parameter GPCFG2_ADDR   = 16'h0008;  //PAD05_CTL  UARTS_TX  0_0001_0000
  parameter GPCFG3_ADDR   = 16'h000C;  //PAD06_CTL  UARTS_RX  0_0000_0111
  parameter GPCFG4_ADDR   = 16'h0010;  //PAD07_CTL  GPIO0     0_0000_0001
  parameter GPCFG5_ADDR   = 16'h0014;  //PAD08_CTL  GPIO1     0_0000_0001
  parameter GPCFG6_ADDR   = 16'h0018;  //PAD09_CTL  GPIO2     0_0000_0001
  parameter GPCFG7_ADDR   = 16'h001C;  //PAD10_CTL  GPIO3     0_0000_0001
  parameter GPCFG8_ADDR   = 16'h0020;  //PAD11_CTL
  parameter GPCFG9_ADDR   = 16'h0024;  //PAD12_CTL
  parameter GPCFG10_ADDR  = 16'h0028;  //PAD13_CTL
  parameter GPCFG11_ADDR  = 16'h002C;  //PAD14_CTL
  parameter GPCFG12_ADDR  = 16'h0030;  //PAD15_CTL
  parameter GPCFG13_ADDR  = 16'h0034;  //PAD16_CTL
  parameter GPCFG14_ADDR  = 16'h0038;  //PAD17_CTL
  parameter GPCFG15_ADDR  = 16'h003C;  //PAD18_CTL
  parameter GPCFG16_ADDR  = 16'h0040;  //PAD19_CTL

  parameter  GPCFG17_ADDR = 16'h0044;  //UARTM_BAUD Reset value for master clock of 25 Mhz and baud rate of 9600
  parameter  GPCFG18_ADDR = 16'h0048;  //UARTM_CTL

  parameter  GPCFG34_ADDR = 16'h0088;  //UARTS_BAUD Reset value for master clock of 25 Mhz and baud rate of 9600
  parameter  GPCFG35_ADDR = 16'h008C;  //UARTS_CTL
  parameter  GPCFG36_ADDR = 16'h0090;  //UARTS_TXDATA
  parameter  GPCFG37_ADDR = 16'h0094;  //UARTS_RXDATA
  parameter  GPCFG38_ADDR = 16'h0098;  //UARTS_TX_SEND
  parameter  GPCFG39_ADDR = 16'h009C;  //SPARE0
  parameter  GPCFG40_ADDR = 16'h00A0;  //SPARE1
  parameter  GPCFG41_ADDR = 16'h00A4;  //SPARE2
  parameter  GPCFG42_ADDR = 16'h00A8;  //CLEEQ_CTL2

  parameter  GPCFG51_ADDR = 16'h00CC;  //SIGNATURE

  parameter  GPCFG_CLCTLP_ADDR      = 16'h8000;
  parameter  GPCFG_CLCTL_ADDR       = 16'h8004;
  parameter  GPCFG_CLSTATUS_ADDR    = 16'h8008;

  parameter [15:0] GPCFG_N_ADDR[0:31] = '{16'h9000,
                                          16'h9004,
                                          16'h9008,
                                          16'h900C,
                                          16'h9010,
                                          16'h9014,
                                          16'h9018,
                                          16'h901C,
                                          16'h9020,
                                          16'h9024,
                                          16'h9028,
                                          16'h902C,
                                          16'h9030,
                                          16'h9034,
                                          16'h9038,
                                          16'h903C,
                                          16'h9040,
                                          16'h9044,
                                          16'h9048,
                                          16'h904C,
                                          16'h9050,
                                          16'h9054,
                                          16'h9058,
                                          16'h905C,
                                          16'h9060,
                                          16'h9064,
                                          16'h9068,
                                          16'h906C,
                                          16'h9070,
                                          16'h9074,
                                          16'h9078,
                                          16'h907C};

  parameter [15:0] GPCFG_R_ADDR[0:31]  = '{16'h9080,
                                           16'h9084,
                                           16'h9088,
                                           16'h908C,
                                           16'h9090,
                                           16'h9094,
                                           16'h9098,
                                           16'h909C,
                                           16'h90A0,
                                           16'h90A4,
                                           16'h90A8,
                                           16'h90AC,
                                           16'h90B0,
                                           16'h90B4,
                                           16'h90B8,
                                           16'h90BC,
                                           16'h90C0,
                                           16'h90C4,
                                           16'h90C8,
                                           16'h90CC,
                                           16'h90D0,
                                           16'h90D4,
                                           16'h90D8,
                                           16'h90DC,
                                           16'h90E0,
                                           16'h90E4,
                                           16'h90E8,
                                           16'h90EC,
                                           16'h90F0,
                                           16'h90F4,
                                           16'h90F8,
                                           16'h90FC};

  parameter [15:0]  GPCFG_NSQ_ADDR[0:63]   = '{16'h9100,
                                               16'h9104,
                                               16'h9108,
                                               16'h910C,
                                               16'h9110,
                                               16'h9114,
                                               16'h9118,
                                               16'h911C,
                                               16'h9120,
                                               16'h9124,
                                               16'h9128,
                                               16'h912C,
                                               16'h9130,
                                               16'h9134,
                                               16'h9138,
                                               16'h913C,
                                               16'h9140,
                                               16'h9144,
                                               16'h9148,
                                               16'h914C,
                                               16'h9150,
                                               16'h9154,
                                               16'h9158,
                                               16'h915C,
                                               16'h9160,
                                               16'h9164,
                                               16'h9168,
                                               16'h916C,
                                               16'h9170,
                                               16'h9174,
                                               16'h9178,
                                               16'h917C,
                                               16'h9180,
                                               16'h9184,
                                               16'h9188,
                                               16'h918C,
                                               16'h9190,
                                               16'h9194,
                                               16'h9198,
                                               16'h919C,
                                               16'h91A0,
                                               16'h91A4,
                                               16'h91A8,
                                               16'h91AC,
                                               16'h91B0,
                                               16'h91B4,
                                               16'h91B8,
                                               16'h91BC,
                                               16'h91C0,
                                               16'h91C4,
                                               16'h91C8,
                                               16'h91CC,
                                               16'h91D0,
                                               16'h91D4,
                                               16'h91D8,
                                               16'h91DC,
                                               16'h91E0,
                                               16'h91E4,
                                               16'h91E8,
                                               16'h91EC,
                                               16'h91F0,
                                               16'h91F4,
                                               16'h91F8,
                                               16'h91FC};

  parameter       [15:0]  GPCFG_FKF_ADDR[0:63]   = '{16'h9200,
                                                     16'h9204,
                                                     16'h9208,
                                                     16'h920C,
                                                     16'h9210,
                                                     16'h9214,
                                                     16'h9218,
                                                     16'h921C,
                                                     16'h9220,
                                                     16'h9224,
                                                     16'h9228,
                                                     16'h922C,
                                                     16'h9230,
                                                     16'h9234,
                                                     16'h9238,
                                                     16'h923C,
                                                     16'h9240,
                                                     16'h9244,
                                                     16'h9248,
                                                     16'h924C,
                                                     16'h9250,
                                                     16'h9254,
                                                     16'h9258,
                                                     16'h925C,
                                                     16'h9260,
                                                     16'h9264,
                                                     16'h9268,
                                                     16'h926C,
                                                     16'h9270,
                                                     16'h9274,
                                                     16'h9278,
                                                     16'h927C,
                                                     16'h9280,
                                                     16'h9284,
                                                     16'h9288,
                                                     16'h928C,
                                                     16'h9290,
                                                     16'h9294,
                                                     16'h9298,
                                                     16'h929C,
                                                     16'h92A0,
                                                     16'h92A4,
                                                     16'h92A8,
                                                     16'h92AC,
                                                     16'h92B0,
                                                     16'h92B4,
                                                     16'h92B8,
                                                     16'h92BC,
                                                     16'h92C0,
                                                     16'h92C4,
                                                     16'h92C8,
                                                     16'h92CC,
                                                     16'h92D0,
                                                     16'h92D4,
                                                     16'h92D8,
                                                     16'h92DC,
                                                     16'h92E0,
                                                     16'h92E4,
                                                     16'h92E8,
                                                     16'h92EC,
                                                     16'h92F0,
                                                     16'h92F4,
                                                     16'h92F8,
                                                     16'h92FC};

  parameter [15:0]  GPCFG_ARGA_ADDR[0:63]   = '{16'h9300,
                                                16'h9304,
                                                16'h9308,
                                                16'h930C,
                                                16'h9310,
                                                16'h9314,
                                                16'h9318,
                                                16'h931C,
                                                16'h9320,
                                                16'h9324,
                                                16'h9328,
                                                16'h932C,
                                                16'h9330,
                                                16'h9334,
                                                16'h9338,
                                                16'h933C,
                                                16'h9340,
                                                16'h9344,
                                                16'h9348,
                                                16'h934C,
                                                16'h9350,
                                                16'h9354,
                                                16'h9358,
                                                16'h935C,
                                                16'h9360,
                                                16'h9364,
                                                16'h9368,
                                                16'h936C,
                                                16'h9370,
                                                16'h9374,
                                                16'h9378,
                                                16'h937C,
                                                16'h9380,
                                                16'h9384,
                                                16'h9388,
                                                16'h938C,
                                                16'h9390,
                                                16'h9394,
                                                16'h9398,
                                                16'h939C,
                                                16'h93A0,
                                                16'h93A4,
                                                16'h93A8,
                                                16'h93AC,
                                                16'h93B0,
                                                16'h93B4,
                                                16'h93B8,
                                                16'h93BC,
                                                16'h93C0,
                                                16'h93C4,
                                                16'h93C8,
                                                16'h93CC,
                                                16'h93D0,
                                                16'h93D4,
                                                16'h93D8,
                                                16'h93DC,
                                                16'h93E0,
                                                16'h93E4,
                                                16'h93E8,
                                                16'h93EC,
                                                16'h93F0,
                                                16'h93F4,
                                                16'h93F8,
                                                16'h93FC};

  parameter [15:0]  GPCFG_ARGB_ADDR[0:63]   = '{16'h9400,
                                                16'h9404,
                                                16'h9408,
                                                16'h940C,
                                                16'h9410,
                                                16'h9414,
                                                16'h9418,
                                                16'h941C,
                                                16'h9420,
                                                16'h9424,
                                                16'h9428,
                                                16'h942C,
                                                16'h9430,
                                                16'h9434,
                                                16'h9438,
                                                16'h943C,
                                                16'h9440,
                                                16'h9444,
                                                16'h9448,
                                                16'h944C,
                                                16'h9450,
                                                16'h9454,
                                                16'h9458,
                                                16'h945C,
                                                16'h9460,
                                                16'h9464,
                                                16'h9468,
                                                16'h946C,
                                                16'h9470,
                                                16'h9474,
                                                16'h9478,
                                                16'h947C,
                                                16'h9480,
                                                16'h9484,
                                                16'h9488,
                                                16'h948C,
                                                16'h9490,
                                                16'h9494,
                                                16'h9498,
                                                16'h949C,
                                                16'h94A0,
                                                16'h94A4,
                                                16'h94A8,
                                                16'h94AC,
                                                16'h94B0,
                                                16'h94B4,
                                                16'h94B8,
                                                16'h94BC,
                                                16'h94C0,
                                                16'h94C4,
                                                16'h94C8,
                                                16'h94CC,
                                                16'h94D0,
                                                16'h94D4,
                                                16'h94D8,
                                                16'h94DC,
                                                16'h94E0,
                                                16'h94E4,
                                                16'h94E8,
                                                16'h94EC,
                                                16'h94F0,
                                                16'h94F4,
                                                16'h94F8,
                                                16'h94FC};

  parameter [15:0]  GPCFG_ARGC_ADDR[0:63]   = '{16'h9500,
                                                16'h9504,
                                                16'h9508,
                                                16'h950C,
                                                16'h9510,
                                                16'h9514,
                                                16'h9518,
                                                16'h951C,
                                                16'h9520,
                                                16'h9524,
                                                16'h9528,
                                                16'h952C,
                                                16'h9530,
                                                16'h9534,
                                                16'h9538,
                                                16'h953C,
                                                16'h9540,
                                                16'h9544,
                                                16'h9548,
                                                16'h954C,
                                                16'h9550,
                                                16'h9554,
                                                16'h9558,
                                                16'h955C,
                                                16'h9560,
                                                16'h9564,
                                                16'h9568,
                                                16'h956C,
                                                16'h9570,
                                                16'h9574,
                                                16'h9578,
                                                16'h957C,
                                                16'h9580,
                                                16'h9584,
                                                16'h9588,
                                                16'h958C,
                                                16'h9590,
                                                16'h9594,
                                                16'h9598,
                                                16'h959C,
                                                16'h95A0,
                                                16'h95A4,
                                                16'h95A8,
                                                16'h95AC,
                                                16'h95B0,
                                                16'h95B4,
                                                16'h95B8,
                                                16'h95BC,
                                                16'h95C0,
                                                16'h95C4,
                                                16'h95C8,
                                                16'h95CC,
                                                16'h95D0,
                                                16'h95D4,
                                                16'h95D8,
                                                16'h95DC,
                                                16'h95E0,
                                                16'h95E4,
                                                16'h95E8,
                                                16'h95EC,
                                                16'h95F0,
                                                16'h95F4,
                                                16'h95F8,
                                                16'h95FC};
  
  parameter [15:0]  GPCFG_RAND0_ADDR[0:31]   = '{16'h9600,
                                                 16'h9604,
                                                 16'h9608,
                                                 16'h960C,
                                                 16'h9610,
                                                 16'h9614,
                                                 16'h9618,
                                                 16'h961C,
                                                 16'h9620,
                                                 16'h9624,
                                                 16'h9628,
                                                 16'h962C,
                                                 16'h9630,
                                                 16'h9634,
                                                 16'h9638,
                                                 16'h963C,
                                                 16'h9640,
                                                 16'h9644,
                                                 16'h9648,
                                                 16'h964C,
                                                 16'h9650,
                                                 16'h9654,
                                                 16'h9658,
                                                 16'h965C,
                                                 16'h9660,
                                                 16'h9664,
                                                 16'h9668,
                                                 16'h966C,
                                                 16'h9670,
                                                 16'h9674,
                                                 16'h9678,
                                                 16'h967C};

  parameter [15:0]  GPCFG_RAND1_ADDR[0:31]       = '{16'h9680,
                                                     16'h9684,
                                                     16'h9688,
                                                     16'h968C,
                                                     16'h9690,
                                                     16'h9694,
                                                     16'h9698,
                                                     16'h969C,
                                                     16'h96A0,
                                                     16'h96A4,
                                                     16'h96A8,
                                                     16'h96AC,
                                                     16'h96B0,
                                                     16'h96B4,
                                                     16'h96B8,
                                                     16'h96BC,
                                                     16'h96C0,
                                                     16'h96C4,
                                                     16'h96C8,
                                                     16'h96CC,
                                                     16'h96D0,
                                                     16'h96D4,
                                                     16'h96D8,
                                                     16'h96DC,
                                                     16'h96E0,
                                                     16'h96E4,
                                                     16'h96E8,
                                                     16'h96EC,
                                                     16'h96F0,
                                                     16'h96F4,
                                                     16'h96F8,
                                                     16'h96FC};

  parameter [15:0]   GPCFG_RES_ADDR[0:63]   = '{16'h9700,
                                                16'h9704,
                                                16'h9708,
                                                16'h970C,
                                                16'h9710,
                                                16'h9714,
                                                16'h9718,
                                                16'h971C,
                                                16'h9720,
                                                16'h9724,
                                                16'h9728,
                                                16'h972C,
                                                16'h9730,
                                                16'h9734,
                                                16'h9738,
                                                16'h973C,
                                                16'h9740,
                                                16'h9744,
                                                16'h9748,
                                                16'h974C,
                                                16'h9750,
                                                16'h9754,
                                                16'h9758,
                                                16'h975C,
                                                16'h9760,
                                                16'h9764,
                                                16'h9768,
                                                16'h976C,
                                                16'h9770,
                                                16'h9774,
                                                16'h9778,
                                                16'h977C,
                                                16'h9780,
                                                16'h9784,
                                                16'h9788,
                                                16'h978C,
                                                16'h9790,
                                                16'h9794,
                                                16'h9798,
                                                16'h979C,
                                                16'h97A0,
                                                16'h97A4,
                                                16'h97A8,
                                                16'h97AC,
                                                16'h97B0,
                                                16'h97B4,
                                                16'h97B8,
                                                16'h97BC,
                                                16'h97C0,
                                                16'h97C4,
                                                16'h97C8,
                                                16'h97CC,
                                                16'h97D0,
                                                16'h97D4,
                                                16'h97D8,
                                                16'h97DC,
                                                16'h97E0,
                                                16'h97E4,
                                                16'h97E8,
                                                16'h97EC,
                                                16'h97F0,
                                                16'h97F4,
                                                16'h97F8,
                                                16'h97FC};

  parameter [15:0]  GPCFG_MUL_ADDR[0:63]   = '{16'h9800,
                                               16'h9804,
                                               16'h9808,
                                               16'h980C,
                                               16'h9810,
                                               16'h9814,
                                               16'h9818,
                                               16'h981C,
                                               16'h9820,
                                               16'h9824,
                                               16'h9828,
                                               16'h982C,
                                               16'h9830,
                                               16'h9834,
                                               16'h9838,
                                               16'h983C,
                                               16'h9840,
                                               16'h9844,
                                               16'h9848,
                                               16'h984C,
                                               16'h9850,
                                               16'h9854,
                                               16'h9858,
                                               16'h985C,
                                               16'h9860,
                                               16'h9864,
                                               16'h9868,
                                               16'h986C,
                                               16'h9870,
                                               16'h9874,
                                               16'h9878,
                                               16'h987C,
                                               16'h9880,
                                               16'h9884,
                                               16'h9888,
                                               16'h988C,
                                               16'h9890,
                                               16'h9894,
                                               16'h9898,
                                               16'h989C,
                                               16'h98A0,
                                               16'h98A4,
                                               16'h98A8,
                                               16'h98AC,
                                               16'h98B0,
                                               16'h98B4,
                                               16'h98B8,
                                               16'h98BC,
                                               16'h98C0,
                                               16'h98C4,
                                               16'h98C8,
                                               16'h98CC,
                                               16'h98D0,
                                               16'h98D4,
                                               16'h98D8,
                                               16'h98DC,
                                               16'h98E0,
                                               16'h98E4,
                                               16'h98E8,
                                               16'h98EC,
                                               16'h98F0,
                                               16'h98F4,
                                               16'h98F8,
                                               16'h98FC};

  parameter [15:0]  GPCFG_EXP_ADDR[0:63]   = '{16'h9900,
                                               16'h9904,
                                               16'h9908,
                                               16'h990C,
                                               16'h9910,
                                               16'h9914,
                                               16'h9918,
                                               16'h991C,
                                               16'h9920,
                                               16'h9924,
                                               16'h9928,
                                               16'h992C,
                                               16'h9930,
                                               16'h9934,
                                               16'h9938,
                                               16'h993C,
                                               16'h9940,
                                               16'h9944,
                                               16'h9948,
                                               16'h994C,
                                               16'h9950,
                                               16'h9954,
                                               16'h9958,
                                               16'h995C,
                                               16'h9960,
                                               16'h9964,
                                               16'h9968,
                                               16'h996C,
                                               16'h9970,
                                               16'h9974,
                                               16'h9978,
                                               16'h997C,
                                               16'h9980,
                                               16'h9984,
                                               16'h9988,
                                               16'h998C,
                                               16'h9990,
                                               16'h9994,
                                               16'h9998,
                                               16'h999C,
                                               16'h99A0,
                                               16'h99A4,
                                               16'h99A8,
                                               16'h99AC,
                                               16'h99B0,
                                               16'h99B4,
                                               16'h99B8,
                                               16'h99BC,
                                               16'h99C0,
                                               16'h99C4,
                                               16'h99C8,
                                               16'h99CC,
                                               16'h99D0,
                                               16'h99D4,
                                               16'h99D8,
                                               16'h99DC,
                                               16'h99E0,
                                               16'h99E4,
                                               16'h99E8,
                                               16'h99EC,
                                               16'h99F0,
                                               16'h99F4,
                                               16'h99F8,
                                               16'h99FC};

  parameter [15:0]  GPCFG_INV_ADDR[0:63]   = '{16'h9A00,
                                               16'h9A04,
                                               16'h9A08,
                                               16'h9A0C,
                                               16'h9A10,
                                               16'h9A14,
                                               16'h9A18,
                                               16'h9A1C,
                                               16'h9A20,
                                               16'h9A24,
                                               16'h9A28,
                                               16'h9A2C,
                                               16'h9A30,
                                               16'h9A34,
                                               16'h9A38,
                                               16'h9A3C,
                                               16'h9A40,
                                               16'h9A44,
                                               16'h9A48,
                                               16'h9A4C,
                                               16'h9A50,
                                               16'h9A54,
                                               16'h9A58,
                                               16'h9A5C,
                                               16'h9A60,
                                               16'h9A64,
                                               16'h9A68,
                                               16'h9A6C,
                                               16'h9A70,
                                               16'h9A74,
                                               16'h9A78,
                                               16'h9A7C,
                                               16'h9A80,
                                               16'h9A84,
                                               16'h9A88,
                                               16'h9A8C,
                                               16'h9A90,
                                               16'h9A94,
                                               16'h9A98,
                                               16'h9A9C,
                                               16'h9AA0,
                                               16'h9AA4,
                                               16'h9AA8,
                                               16'h9AAC,
                                               16'h9AB0,
                                               16'h9AB4,
                                               16'h9AB8,
                                               16'h9ABC,
                                               16'h9AC0,
                                               16'h9AC4,
                                               16'h9AC8,
                                               16'h9ACC,
                                               16'h9AD0,
                                               16'h9AD4,
                                               16'h9AD8,
                                               16'h9ADC,
                                               16'h9AE0,
                                               16'h9AE4,
                                               16'h9AE8,
                                               16'h9AEC,
                                               16'h9AF0,
                                               16'h9AF4,
                                               16'h9AF8,
                                               16'h9AFC};


  parameter [15:0]  GPCFG_DBG_ADDR[0:63]   = '{16'h9B00,
                                               16'h9B04,
                                               16'h9B08,
                                               16'h9B0C,
                                               16'h9B10,
                                               16'h9B14,
                                               16'h9B18,
                                               16'h9B1C,
                                               16'h9B20,
                                               16'h9B24,
                                               16'h9B28,
                                               16'h9B2C,
                                               16'h9B30,
                                               16'h9B34,
                                               16'h9B38,
                                               16'h9B3C,
                                               16'h9B40,
                                               16'h9B44,
                                               16'h9B48,
                                               16'h9B4C,
                                               16'h9B50,
                                               16'h9B54,
                                               16'h9B58,
                                               16'h9B5C,
                                               16'h9B60,
                                               16'h9B64,
                                               16'h9B68,
                                               16'h9B6C,
                                               16'h9B70,
                                               16'h9B74,
                                               16'h9B78,
                                               16'h9B7C,
                                               16'h9B80,
                                               16'h9B84,
                                               16'h9B88,
                                               16'h9B8C,
                                               16'h9B90,
                                               16'h9B94,
                                               16'h9B98,
                                               16'h9B9C,
                                               16'h9BA0,
                                               16'h9BA4,
                                               16'h9BA8,
                                               16'h9BAC,
                                               16'h9BB0,
                                               16'h9BB4,
                                               16'h9BB8,
                                               16'h9BBC,
                                               16'h9BC0,
                                               16'h9BC4,
                                               16'h9BC8,
                                               16'h9BCC,
                                               16'h9BD0,
                                               16'h9BD4,
                                               16'h9BD8,
                                               16'h9BDC,
                                               16'h9BE0,
                                               16'h9BE4,
                                               16'h9BE8,
                                               16'h9BEC,
                                               16'h9BF0,
                                               16'h9BF4,
                                               16'h9BF8,
                                               16'h9BFC};


